module mul32p_tb(
    
);
endmodule