module mul_tb_qhw;
endmodule